b0VIM 8.2      �l�f " root                                    vps-9ecac94e                            /var/www/veopro/VEO/models.py                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           �                     ��������_       �              ��������O       �              ��������F       1             ��������]       w             ��������Q       �             ��������_       %             ��������K       �             ��������6       �             ��������P                    ��������^       U             ��������6       �             ��������R       �             ��������@       ;             ��������M       {             ��������N       �             ��������1                    ��������1       G                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ad     B     �       �  �  �  �  �    m    �  �  �  �  �  �  �  s  c  b  a  `  _  D  )    �  �  }  c  K    �  �  �  Y  ;      �  �  �  �  �  �  �  p  ^  E  #    �
  �
  �
  �
  �
  �
  |
  i
  M
  .
  
  �	  �	  �	  �	  �	  �	  �	  	  [	  P	  ?	  >	  =	  	  �  �  �  j  N  0      �  �  �  �  �  y  N    �  �  �  �  �  �  s  X  H  0      �  �  �  �  x  Z  C  +    �  w  `  K  J  '  �  �  �  �  }  e  d  G    �  �  i  B  A                                    Immatriculation=models.TextField()     ContactName=models.TextField()     Type=models.TextField()     Collaborateur = models.ForeignKey(Collaborateur, on_delete=models.SET_NULL, null=True, related_name='veodata')     id = models.TextField(primary_key=True) class Veodata(models.Model):          return self.nom     def __str__(self):      nom = models.TextField(max_length=100)     email = models.EmailField(max_length=254, unique=True)     id = models.TextField(primary_key=True) class Collaborateur(models.Model):              return a             #a=test(a)             # cette fonction élimine les immatriculation qui sont tous des zéros et qui sont tous des lettres              a=add_zero(a)         if (a != '' and not(a is None)):         a=remove_WW0(a)         a=remove_WW(a)         a=remove_zerostart(a)         a=a.replace('-','')         a=a.replace(".", "")         a=a.replace("'", "")         a=a.replace("/", "")         a=a.replace(" ", "")         a=a.upper()         a=a.strip()         a=remove_EAD(a)     if a!=None: def Preprocessing_Imm (a): #Preprocessing "Immatriculation" (Appeler toutes les fcts défénies)           return a     else:         return ""     if ((len(b) == len(a)) or ((len(c) == len(a)))):     c=''.join(i for i in a if not (i.isdigit()))     b=''.join(i for i in a if i.isdigit()) def test(a): #Enlever les imm qui contient que des chiffres ou bien que des caractères          return a     else:             return a         else:             return ''.join(res)             res.append(a[-1])             res.append("0")             res=list(a)[0:-1]         if (a[-1].isdigit() and (not a[-2].isdigit())):     if (len(a) <= 2 or a != '' or not (a is None)): def add_zero(a): #Ajouter le le zéro après le caractère (B7 ==> B07)            return a     else:          return ''.join(list(a)[3:])     if (a.startswith("EAD")): def remove_EAD(a): #Enlever le mot "EAD" s'il existe          return a     else:         return a         a="WW"+a         a=remove_zerostart(a)         a=''.join(list(a)[2:])     if a.startswith("WW0"): def remove_WW0(a): #Enlever les zeros après les "WW" de début          return a     else:             return "WW"+a         else :             return a         if(a.startswith("WW")):         a= ''.join(list(a)[0:-2])     if a.endswith("WW"): def remove_WW(a): #Enlever les "WW" à la fin      return val         val = ''.join(l)         i=i+1         l[0]=''         l=list(val)     while (val.startswith('0') and i<len(val)):     i=0 def remove_zerostart (val): #Enlever les zéros de début ############################################################### Nettoyage des immatriculations          return abs(dtE- dtV).days          dtE = datetime.strptime(dtE, "%d/%m/%Y").date()         dtV= datetime.strptime(dtV, "%d/%m/%Y").date()     if (dtV and dtE):   def inter_dt2(dtV,dtE):           return abs(dtV - dtE).days          dtE = datetime.strptime(dtE, "%d/%m/%Y").date()         dtV = datetime.strptime(dtV, "%d/%m/%Y").date()     if (dtV and dtE):   def inter_dt(dtV , dtE):   # Create your models here.         return stri         stri=float(stri)     else:         stri=0.0     if stri == "" or stri == "'0.0'" or stri  == None: def str_to_float(stri):       return a     a=a.replace(' ','').replace('-','').replace('_','').replace(',','').replace('.','').replace('*','') def net_numch(a): # nettoyage  de  numéro de  chassis   from django.db.models import Q from datetime import datetime from django.db import models ad  J  *     1       �  �  2      �  �  �  N  7  6         �
  j
  ]
  q	  p	  X	  �  �  �  x  w  _  �  �  �  �  y  Z  Y  X  C  4  %  �  �  �  ]  I  H  ?  :  9  8  /  *  )                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   return Rate         veotest.objects.filter(id=self.id).update(R14=R)              R="Ce sinistre est en instruction"             Rate=15         if (self.statutdt_omega == "Dossier initié" or self.statutdt_omega == "Dossier initié RMAA" or self.statutdt_omega == "Doute créé" or self.statutdt_omega == "Dossier envoyé"  or self.statutdt_omega == "Affecté expert" or self.statutdt_omega == "Retour expert" or self.statutdt_omega == "Attente photos avant")  :             Rate=0         R=None     def Reg14(self):               return [Rate,Doss]             veotest.objects.filter(id=self.id).update(R13=R)                                Doss=i                 R="l'immatriculation Adverse a déjà été impliquée dans un dossier historique doute rejeté : "+str(i.Dossier)                 Rate=15              elif i.Immatriculation != "" and self.Immatriculation != "" and i.ImmatriculationAdverse != "" and self.ImmatriculationAdverse != "" and i.ImmatriculationAdverse == self.ImmatriculationAdverse and (i.statutdt_omega != "Doute rejeté" or i.statutdt_omega != "Doute rejeté RMAA")  and i.statutdt_omega != None:                  Doss=i                 R="l'immatriculation principale a déjà été impliquée dans un dossier historique doute rejeté : "+str(i.Dossier)                 Rate=15              elif i.Immatriculation != "" and self.Immatriculation != ""  and i.Immatriculation == self.Immatriculation and (i.statutdt_omega != "Doute rejeté" or i.statutdt_omega != "Doute rejeté RMAA")  and i.statutdt_omega != None:                              Doss=i                 R="l'immatriculation principale a déjà été impliquée dans un dossier historique doute rejeté : "+str(i.Dossier)                 Rate=15              elif i.Immatriculation != "" and self.Immatriculation != "" and i.ImmatriculationAdverse != ""  and i.ImmatriculationAdverse == self.Immatriculation and (i.statutdt_omega != "Doute rejeté" or i.statutdt_omega != "Doute rejeté RMAA")  and i.statutdt_omega != None:                  Doss=i                 R="l'immatriculation Adverse a déjà été impliquée dans un dossier historique doute rejeté : "+str(i.Dossier)                 Rate=15              elif i.Immatriculation != "" and self.Immatriculation != ""  and  self.ImmatriculationAdverse != ""  and i.Immatriculation == self.ImmatriculationAdverse and (i.statutdt_omega != "Doute rejeté" or i.statutdt_omega != "Doute rejeté RMAA")  and i.statutdt_omega != None:                                       Doss=i                 R="l'immatriculation Adverse a déjà été impliquée dans un dossier historique doute confirmé : "+str(i.Dossier)                 Rate=30             elif i.Immatriculation != "" and self.Immatriculation != ""  and i.ImmatriculationAdverse != "" and self.ImmatriculationAdverse != ""  and i.ImmatriculationAdverse == self.ImmatriculationAdverse and (i.statutdt_omega == "Doute confirmé" or i.statutdt_omega == "Doute confirmé RMAA" )  :     